`define ON_1b 1'b1
`define OFF_1b 1'b0
`define UNPLUGED 1'bz
`define NM_1b 1'bx

`define ON_2b 2'b1
`define OFF_2b 2'b0

`define ON_3b 3'b1
`define OFF_3b 3'b0 