`define MIPS_ADD   6'h20
`define MIPS_SUB   6'h22
`define MIPS_AND   6'h24
`define MIPS_OR    6'h25
`define MIPS_SLT   6'h2A
`define MIPS_LW    6'h23
`define MIPS_SW    6'h2B
`define MIPS_BEQ   6'h04
`define MIPS_BNE   6'h05
`define MIPS_JUMP  6'h02

`define MIPS_ADDU  6'h21
`define MIPS_SUBU  6'h23
`define MIPS_ADDI  6'h08
`define MIPS_ADDIU 6'h09
`define MIPS_ANDI  6'h0C
`define MIPS_ORI   6'h0D
`define MIPS_LUI   6'h0F
`define MIPS_XOR   6'h26
`define MIPS_XORI  6'h0E
`define MIPS_SLTI  6'h0A
`define MIPS_SLTU  6'h2B
`define MIPS_SLTIU 6'h0B

`define MIPS_LH    6'h21
`define MIPS_LHU   6'h25
`define MIPS_LB    6'h20
`define MIPS_LBU   6'h24
`define MIPS_SH    6'h29
`define MIPS_SB    6'h28

